module gates_using_nand_tb;
	// Inputs
	reg a;
	reg b;
	// Outputs
	wire y;

	// Instantiate the Unit Under Test (UUT)
	gates_using_nand uut (.a(a), .b(b), .y(y));

	initial begin
		// Initialize Inputs
		a = 0;
		b = 0;
		#10;        
		// Add stimulus here
		a = 0;
		b = 1;
		#10; 
		a = 1;
		b = 0;
		#10;       
		a = 1;
		b = 1;
		#10;      		 
	end
	initial 
		begin
			$monitor("a=%b,b=%b,y=%b",a,b,y);
		end      
endmodule
