module jk_latch (
  input j,
  input k,
  input en,        // enable or clock input
  output reg q,
  output qbar
);
  assign qbar = ~q;

  always @(*) begin
    if (en) begin
      case ({j, k})
        2'b00: q = q;      // Hold
        2'b01: q = 1'b0;   // Reset
        2'b10: q = 1'b1;   // Set
        2'b11: q = ~q;     // Toggle
      endcase
    end
  end
endmodule
